----------------------------------------------------------------------------------
------------------------------EXPANSION-PERMUTATION-BOX---------------------------
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


--entity
entity EXP_BOX is
    port(STD_LOGIC_1164
        INPUT: IN STD_LOGIC_VECTOR(31 downto 0);
        OUTPUT: OUT STD_LOGIC_VECTOR(47 downto 0)
    )
end EXP_BOX;


--architecture
architecture Behavioral of EXP_BOX is

begin


end Behavioral;

